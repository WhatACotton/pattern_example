/* Copyright(C) 2020 Cobac.Net All Rights Reserved. */
/* chapter: 第2章                     */
/* project: pattern                   */
/* outline: ピクセルクロック生成      */
/*          125MHz入力、25.175MHz出力 */

`ifndef SYNTHESIS
`include "../imports/src/rgb2dvi.vhd"
`endif
module pckgen (
    input  SYSCLK,
    output PCK
);

  wire CLKFBOUT, iPCK, locked;
  BUFG iBUFG (
      .I(iPCK),
      .O(PCK)
  );

  MMCME2_BASE #(
      .BANDWIDTH         ("OPTIMIZED"),  // Jitter programming (OPTIMIZED, HIGH, LOW)
      .CLKFBOUT_MULT_F   (36.0),         // 乗数M(2.000-64.000)
      .CLKFBOUT_PHASE    (0.0),          // 位相(-360.000-360.000)
      .CLKIN1_PERIOD     (8.0),          // CLKINの周期
      // CLKOUT0_DIVIDE - CLKOUT6_DIVIDE: Divide amount for each CLKOUT (1-128)
      .CLKOUT1_DIVIDE    (1),
      .CLKOUT2_DIVIDE    (1),
      .CLKOUT3_DIVIDE    (1),
      .CLKOUT4_DIVIDE    (1),
      .CLKOUT5_DIVIDE    (1),
      .CLKOUT6_DIVIDE    (1),
      .CLKOUT0_DIVIDE_F  (35.75),        // 除数Q(1.000-128.000)
      // CLKOUT0_DUTY_CYCLE - CLKOUT6_DUTY_CYCLE: Duty cycle for each CLKOUT (0.01-0.99).
      .CLKOUT0_DUTY_CYCLE(0.5),          // デューティ比
      .CLKOUT1_DUTY_CYCLE(0.5),
      .CLKOUT2_DUTY_CYCLE(0.5),
      .CLKOUT3_DUTY_CYCLE(0.5),
      .CLKOUT4_DUTY_CYCLE(0.5),
      .CLKOUT5_DUTY_CYCLE(0.5),
      .CLKOUT6_DUTY_CYCLE(0.5),
      // CLKOUT0_PHASE - CLKOUT6_PHASE: Phase offset for each CLKOUT (-360.000-360.000).
      .CLKOUT0_PHASE     (0.0),
      .CLKOUT1_PHASE     (0.0),
      .CLKOUT2_PHASE     (0.0),
      .CLKOUT3_PHASE     (0.0),
      .CLKOUT4_PHASE     (0.0),
      .CLKOUT5_PHASE     (0.0),
      .CLKOUT6_PHASE     (0.0),
      .CLKOUT4_CASCADE   ("FALSE"),      // Cascade CLKOUT4 counter with CLKOUT6 (FALSE, TRUE)
      .DIVCLK_DIVIDE     (5),            // 除数D(1-106)
      .REF_JITTER1       (0.0),          // Reference input jitter in UI (0.000-0.999).
      .STARTUP_WAIT      ("FALSE")       // Delays DONE until MMCM is locked (FALSE, TRUE)
  ) MMCME2_BASE_inst (
      // Clock Outputs: 1-bit (each) output: User configurable clock outputs
      .CLKOUT0  (iPCK),      // 1-bit output: CLKOUT0
      .CLKOUT0B (),          // 1-bit output: Inverted CLKOUT0
      .CLKOUT1  (),          // 1-bit output: CLKOUT1
      .CLKOUT1B (),          // 1-bit output: Inverted CLKOUT1
      .CLKOUT2  (),          // 1-bit output: CLKOUT2
      .CLKOUT2B (),          // 1-bit output: Inverted CLKOUT2
      .CLKOUT3  (),          // 1-bit output: CLKOUT3
      .CLKOUT3B (),          // 1-bit output: Inverted CLKOUT3
      .CLKOUT4  (),          // 1-bit output: CLKOUT4
      .CLKOUT5  (),          // 1-bit output: CLKOUT5
      .CLKOUT6  (),          // 1-bit output: CLKOUT6
      // Feedback Clocks: 1-bit (each) output: Clock feedback ports
      .CLKFBOUT (CLKFBOUT),  // 1-bit output: Feedback clock
      .CLKFBOUTB(),          // 1-bit output: Inverted CLKFBOUT
      // Status Ports: 1-bit (each) output: MMCM status ports
      .LOCKED   (locked),    // 1-bit output: LOCK
      // Clock Inputs: 1-bit (each) input: Clock input
      .CLKIN1   (SYSCLK),    // 1-bit input: Clock
      // Control Ports: 1-bit (each) input: MMCM control ports
      .PWRDWN   (1'b0),      // 1-bit input: Power-down
      .RST      (1'b0),      // 1-bit input: Reset
      // Feedback Clocks: 1-bit (each) input: Clock feedback ports
      .CLKFBIN  (CLKFBOUT)   // 1-bit input: Feedback clock
  );

endmodule
